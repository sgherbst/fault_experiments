`timescale 1ns/1ns
module sram_2_16_scn4m_subm_tb;
    reg [1:0] din0;
    wire [1:0] dout0;
    reg [3:0] addr0;
    reg csb0;
    reg web0;
    reg clk0;

    

    sram_2_16_scn4m_subm #(
        
    ) dut (
        .din0(din0),
        .dout0(dout0),
        .addr0(addr0),
        .csb0(csb0),
        .web0(web0),
        .clk0(clk0)
    );

    initial begin
        $dumpfile("waveforms.vcd");
        $dumpvars(0, dut);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        csb0 <= 1'b0;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(5e-08*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(5e-08*1s);
        din0 <= 2'd1;
        #(0*1s);
        addr0 <= 4'd3;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd6;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd8;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd1;
        #(0*1s);
        addr0 <= 4'd2;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd5;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd12;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd15;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd11;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd14;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd4;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd1;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd13;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd10;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd9;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd7;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        addr0 <= 4'd6;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=193 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=203 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd7;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=213 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd10;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=223 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd3;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd1)) begin
            $error("Failed on action=233 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd1, dout0);
        end
        addr0 <= 4'd12;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=243 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd14;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=253 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd11;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=263 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd9;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=273 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd15;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=283 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd4;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=293 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd1;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=303 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd8;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=313 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd13;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=323 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd5;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=333 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd2;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd1)) begin
            $error("Failed on action=343 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd1, dout0);
        end
        #20 $finish;
    end

endmodule

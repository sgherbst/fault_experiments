* Automatically generated file.
.include /Users/sgherbst/Dropbox/LaptopSync/Stanford/Research/Code/fault_experiments/sram/nmos.sp
.include /Users/sgherbst/Dropbox/LaptopSync/Stanford/Research/Code/fault_experiments/sram/pmos.sp
.include /Users/sgherbst/Dropbox/LaptopSync/Stanford/Research/Code/fault_experiments/sram/sram_8_16_scn4m_subm.sp
X0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] addr0[0] addr0[1] addr0[2] addr0[3] csb0 web0 clk0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] vdd gnd sram_8_16_scn4m_subm
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    Gs sw_p sw_n cur='V(sw_p, sw_n)*(0.999999999*V(ctl_p, ctl_n)+1e-09)'
.ends
X1 __din0[0]_v din0[0] __din0[0]_s 0 inout_sw_mod
V2 __din0[0]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 0 5.6e-08 0 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 0 1.0599999999999998e-07 0 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 0 1.1599999999999998e-07 0 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V3 __din0[0]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X4 __din0[1]_v din0[1] __din0[1]_s 0 inout_sw_mod
V5 __din0[1]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 0 7.599999999999999e-08 0 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 0 1.1599999999999998e-07 0 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V6 __din0[1]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X7 __din0[2]_v din0[2] __din0[2]_s 0 inout_sw_mod
V8 __din0[2]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 3.3 6.6e-08 3.3 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 3.3 8.599999999999999e-08 3.3 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 3.3 9.599999999999999e-08 3.3 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V9 __din0[2]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X10 __din0[3]_v din0[3] __din0[3]_s 0 inout_sw_mod
V11 __din0[3]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 3.3 6.6e-08 3.3 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 3.3 8.599999999999999e-08 3.3 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 0 1.0599999999999998e-07 0 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V12 __din0[3]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X13 __din0[4]_v din0[4] __din0[4]_s 0 inout_sw_mod
V14 __din0[4]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 0 5.6e-08 0 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 0 7.599999999999999e-08 0 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 3.3 9.599999999999999e-08 3.3 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V15 __din0[4]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X16 __din0[5]_v din0[5] __din0[5]_s 0 inout_sw_mod
V17 __din0[5]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 3.3 6.6e-08 3.3 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 0 1.1599999999999998e-07 0 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V18 __din0[5]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X19 __din0[6]_v din0[6] __din0[6]_s 0 inout_sw_mod
V20 __din0[6]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 3.3 8.599999999999999e-08 3.3 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 0 1.1599999999999998e-07 0 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V21 __din0[6]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X22 __din0[7]_v din0[7] __din0[7]_s 0 inout_sw_mod
V23 __din0[7]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 3.3 6.6e-08 3.3 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 3.3 9.599999999999999e-08 3.3 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 3.700000000000002e-07 0)
V24 __din0[7]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 3.700000000000002e-07 1)
X25 __addr0[0]_v addr0[0] __addr0[0]_s 0 inout_sw_mod
V26 __addr0[0]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 0 5.6e-08 0 5.62e-08 0 6e-08 0 6.02e-08 3.3 6.6e-08 3.3 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 0 7.599999999999999e-08 0 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 3.3 9.599999999999999e-08 3.3 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 0 1.46e-07 0 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 0 2.6600000000000013e-07 0 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 0 2.7600000000000014e-07 0 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 0 2.8600000000000015e-07 0 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 0 3.0600000000000017e-07 0 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 0 3.160000000000002e-07 0 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 0 3.460000000000002e-07 0 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 3.3 3.560000000000002e-07 3.3 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.700000000000002e-07 0)
V27 __addr0[0]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1)
X28 __addr0[1]_v addr0[1] __addr0[1]_s 0 inout_sw_mod
V29 __addr0[1]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 0 5.6e-08 0 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 3.3 9.599999999999999e-08 3.3 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 0 2.6600000000000013e-07 0 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 0 2.8600000000000015e-07 0 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 0 3.260000000000002e-07 0 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 0 3.360000000000002e-07 0 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 0 3.560000000000002e-07 0 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.700000000000002e-07 0)
V30 __addr0[1]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1)
X31 __addr0[2]_v addr0[2] __addr0[2]_s 0 inout_sw_mod
V32 __addr0[2]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 3.3 8.599999999999999e-08 3.3 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 0 1.1599999999999998e-07 0 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 0 2.7600000000000014e-07 0 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 0 3.160000000000002e-07 0 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 0 3.260000000000002e-07 0 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 0 3.560000000000002e-07 0 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 0 3.6600000000000023e-07 0 3.6620000000000025e-07 0 3.700000000000002e-07 0)
V33 __addr0[2]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1)
X34 __addr0[3]_v addr0[3] __addr0[3]_s 0 inout_sw_mod
V35 __addr0[3]_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 5.6e-08 3.3 5.62e-08 0 6e-08 0 6.02e-08 0 6.6e-08 0 6.62e-08 0 6.999999999999999e-08 0 7.019999999999999e-08 0 7.599999999999999e-08 0 7.62e-08 0 7.999999999999999e-08 0 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 0 8.999999999999999e-08 0 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 0 9.999999999999998e-08 0 1.0019999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.0999999999999998e-07 0 1.1019999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 0 2.6600000000000013e-07 0 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 0 2.9600000000000016e-07 0 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 0 3.0600000000000017e-07 0 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 0 3.160000000000002e-07 0 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 0 3.260000000000002e-07 0 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 3.3 3.560000000000002e-07 3.3 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.700000000000002e-07 0)
V36 __addr0[3]_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1)
X37 __csb0_v csb0 __csb0_s 0 inout_sw_mod
V38 __csb0_v 0 DC 0 PWL(0 0 3.700000000000002e-07 0)
V39 __csb0_s 0 DC 1 PWL(0 1 3.700000000000002e-07 1)
X40 __web0_v web0 __web0_s 0 inout_sw_mod
V41 __web0_v 0 DC 0 PWL(0 0 2.5e-08 0 2.5199999999999997e-08 3.3 5e-08 3.3 5.02e-08 0 5.6e-08 0 5.62e-08 3.3 6e-08 3.3 6.02e-08 0 6.6e-08 0 6.62e-08 3.3 6.999999999999999e-08 3.3 7.019999999999999e-08 0 7.599999999999999e-08 0 7.62e-08 3.3 7.999999999999999e-08 3.3 8.019999999999999e-08 0 8.599999999999999e-08 0 8.619999999999999e-08 3.3 8.999999999999999e-08 3.3 9.019999999999999e-08 0 9.599999999999999e-08 0 9.619999999999999e-08 3.3 9.999999999999998e-08 3.3 1.0019999999999998e-07 0 1.0599999999999998e-07 0 1.0619999999999998e-07 3.3 1.0999999999999998e-07 3.3 1.1019999999999998e-07 0 1.1599999999999998e-07 0 1.1619999999999998e-07 3.3 1.2e-07 3.3 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 3.3 1.3e-07 3.3 1.302e-07 0 1.36e-07 0 1.362e-07 3.3 1.4e-07 3.3 1.402e-07 0 1.46e-07 0 1.462e-07 3.3 1.5000000000000002e-07 3.3 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 3.3 1.6000000000000003e-07 3.3 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 3.3 1.7000000000000004e-07 3.3 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 3.3 1.8000000000000005e-07 3.3 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 3.3 1.9000000000000006e-07 3.3 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 3.3 2.0000000000000007e-07 3.3 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 3.3 2.1000000000000008e-07 3.3 2.1020000000000007e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 3.3 2.200000000000001e-07 3.3 2.2020000000000008e-07 3.3 2.260000000000001e-07 3.3 2.2620000000000008e-07 3.3 2.300000000000001e-07 3.3 2.302000000000001e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 3.3 2.400000000000001e-07 3.3 2.402000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 3.3 2.500000000000001e-07 3.3 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 3.3 2.600000000000001e-07 3.3 2.602000000000001e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 3.3 2.700000000000001e-07 3.3 2.7020000000000013e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 3.3 2.800000000000001e-07 3.3 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 3.3 2.9000000000000014e-07 3.3 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 3.3 3.0000000000000015e-07 3.3 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 3.3 3.1000000000000016e-07 3.3 3.1020000000000017e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 3.3 3.2000000000000017e-07 3.3 3.202000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 3.3 3.300000000000002e-07 3.3 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 3.3 3.400000000000002e-07 3.3 3.402000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 3.3 3.500000000000002e-07 3.3 3.502000000000002e-07 3.3 3.560000000000002e-07 3.3 3.5620000000000024e-07 3.3 3.600000000000002e-07 3.3 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 3.3 3.700000000000002e-07 3.3)
V42 __web0_s 0 DC 1 PWL(0 1 2.5e-08 1 2.5199999999999997e-08 1 5e-08 1 5.02e-08 1 5.6e-08 1 5.62e-08 1 6e-08 1 6.02e-08 1 6.6e-08 1 6.62e-08 1 6.999999999999999e-08 1 7.019999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 7.999999999999999e-08 1 8.019999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 8.999999999999999e-08 1 9.019999999999999e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 9.999999999999998e-08 1 1.0019999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.0999999999999998e-07 1 1.1019999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1)
X43 __clk0_v clk0 __clk0_s 0 inout_sw_mod
V44 __clk0_v 0 DC 0 PWL(0 0 5.1e-08 0 5.12e-08 3.3 5.6e-08 3.3 5.62e-08 0 6.099999999999999e-08 0 6.119999999999999e-08 3.3 6.6e-08 3.3 6.62e-08 0 7.099999999999999e-08 0 7.119999999999999e-08 3.3 7.599999999999999e-08 3.3 7.62e-08 0 8.099999999999998e-08 0 8.119999999999999e-08 3.3 8.599999999999999e-08 3.3 8.619999999999999e-08 0 9.099999999999998e-08 0 9.119999999999998e-08 3.3 9.599999999999999e-08 3.3 9.619999999999999e-08 0 1.0099999999999998e-07 0 1.0119999999999998e-07 3.3 1.0599999999999998e-07 3.3 1.0619999999999998e-07 0 1.1099999999999997e-07 0 1.1119999999999998e-07 3.3 1.1599999999999998e-07 3.3 1.1619999999999998e-07 0 1.2099999999999998e-07 0 1.2119999999999997e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.31e-07 0 1.3119999999999998e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.41e-07 0 1.412e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5100000000000002e-07 0 1.512e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6100000000000003e-07 0 1.6120000000000001e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7100000000000004e-07 0 1.7120000000000002e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8100000000000005e-07 0 1.8120000000000003e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9100000000000006e-07 0 1.9120000000000004e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0100000000000007e-07 0 2.0120000000000005e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1100000000000008e-07 0 2.1120000000000006e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 0 2.2100000000000009e-07 0 2.2120000000000007e-07 3.3 2.260000000000001e-07 3.3 2.2620000000000008e-07 0 2.310000000000001e-07 0 2.3120000000000009e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 0 2.410000000000001e-07 0 2.412000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 0 2.510000000000001e-07 0 2.5120000000000013e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.6100000000000013e-07 0 2.6120000000000014e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 0 2.7100000000000014e-07 0 2.7120000000000015e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 0 2.8100000000000015e-07 0 2.8120000000000016e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9100000000000016e-07 0 2.9120000000000017e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0100000000000017e-07 0 3.012000000000002e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.110000000000002e-07 0 3.112000000000002e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 0 3.210000000000002e-07 0 3.212000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 0 3.310000000000002e-07 0 3.312000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.410000000000002e-07 0 3.412000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 0 3.510000000000002e-07 0 3.5120000000000023e-07 3.3 3.560000000000002e-07 3.3 3.5620000000000024e-07 0 3.6100000000000023e-07 0 3.6120000000000024e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.700000000000002e-07 0)
V45 __clk0_s 0 DC 1 PWL(0 1 5.1e-08 1 5.12e-08 1 5.6e-08 1 5.62e-08 1 6.099999999999999e-08 1 6.119999999999999e-08 1 6.6e-08 1 6.62e-08 1 7.099999999999999e-08 1 7.119999999999999e-08 1 7.599999999999999e-08 1 7.62e-08 1 8.099999999999998e-08 1 8.119999999999999e-08 1 8.599999999999999e-08 1 8.619999999999999e-08 1 9.099999999999998e-08 1 9.119999999999998e-08 1 9.599999999999999e-08 1 9.619999999999999e-08 1 1.0099999999999998e-07 1 1.0119999999999998e-07 1 1.0599999999999998e-07 1 1.0619999999999998e-07 1 1.1099999999999997e-07 1 1.1119999999999998e-07 1 1.1599999999999998e-07 1 1.1619999999999998e-07 1 1.2099999999999998e-07 1 1.2119999999999997e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.31e-07 1 1.3119999999999998e-07 1 1.36e-07 1 1.362e-07 1 1.41e-07 1 1.412e-07 1 1.46e-07 1 1.462e-07 1 1.5100000000000002e-07 1 1.512e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6100000000000003e-07 1 1.6120000000000001e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7100000000000004e-07 1 1.7120000000000002e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8100000000000005e-07 1 1.8120000000000003e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9100000000000006e-07 1 1.9120000000000004e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0100000000000007e-07 1 2.0120000000000005e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1100000000000008e-07 1 2.1120000000000006e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.2100000000000009e-07 1 2.2120000000000007e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.310000000000001e-07 1 2.3120000000000009e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.410000000000001e-07 1 2.412000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.510000000000001e-07 1 2.5120000000000013e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.6100000000000013e-07 1 2.6120000000000014e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.7100000000000014e-07 1 2.7120000000000015e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.8100000000000015e-07 1 2.8120000000000016e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9100000000000016e-07 1 2.9120000000000017e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0100000000000017e-07 1 3.012000000000002e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.110000000000002e-07 1 3.112000000000002e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.210000000000002e-07 1 3.212000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.310000000000002e-07 1 3.312000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.410000000000002e-07 1 3.412000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.510000000000002e-07 1 3.5120000000000023e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.6100000000000023e-07 1 3.6120000000000024e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1)
X46 __vdd_v vdd __vdd_s 0 inout_sw_mod
V47 __vdd_v 0 DC 0 PWL(0 0 2.5e-08 0 2.5199999999999997e-08 3.3 3.700000000000002e-07 3.3)
V48 __vdd_s 0 DC 1 PWL(0 1 2.5e-08 1 2.5199999999999997e-08 1 3.700000000000002e-07 1)
X49 __gnd_v gnd __gnd_s 0 inout_sw_mod
V50 __gnd_v 0 DC 0 PWL(0 0 3.700000000000002e-07 0)
V51 __gnd_s 0 DC 1 PWL(0 1 3.700000000000002e-07 1)
.tran 3.700000000000002e-10 3.700000000000002e-07 uic
.control
run
set filetype=binary
write
exit
.endc
.probe V(addr0[3]) V(clk0) V(dout0[7]) V(addr0[0]) V(din0[5]) V(dout0[3]) V(din0[7]) V(din0[0]) V(din0[2]) V(dout0[1]) V(web0) V(vdd) V(gnd) V(din0[1]) V(dout0[6]) V(dout0[2]) V(din0[6]) V(dout0[0]) V(csb0) V(din0[4]) V(addr0[2]) V(din0[3]) V(dout0[4]) V(dout0[5]) V(addr0[1])
.end

`timescale 1ns/1ns
module sram_2_16_scn4m_subm_tb;
    reg [1:0] din0;
    wire [1:0] __din0_wire;
    wire [1:0] dout0;
    reg [3:0] addr0;
    wire [3:0] __addr0_wire;
    reg csb0;
    wire __csb0_wire;
    reg web0;
    wire __web0_wire;
    reg clk0;
    wire __clk0_wire;
    reg vdd;
    wire __vdd_wire;
    reg gnd;
    wire __gnd_wire;
    assign __din0_wire=din0;
    assign __addr0_wire=addr0;
    assign __csb0_wire=csb0;
    assign __web0_wire=web0;
    assign __clk0_wire=clk0;
    assign __vdd_wire=vdd;
    assign __gnd_wire=gnd;
    

    sram_2_16_scn4m_subm #(
        
    ) dut (
        .din0(__din0_wire),
        .dout0(dout0),
        .addr0(__addr0_wire),
        .csb0(__csb0_wire),
        .web0(__web0_wire),
        .clk0(__clk0_wire),
        .vdd(__vdd_wire),
        .gnd(__gnd_wire)
    );

    initial begin
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        csb0 <= 1'b0;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        vdd <= 1'b0;
        #(0*1s);
        gnd <= 1'b0;
        #(0*1s);
        #(5e-08*1s);
        vdd <= 1'b1;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(5e-08*1s);
        din0 <= 2'd1;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd11;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd13;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd9;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd15;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd14;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd8;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd3;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd1;
        #(0*1s);
        addr0 <= 4'd2;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd5;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd1;
        #(0*1s);
        addr0 <= 4'd12;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd3;
        #(0*1s);
        addr0 <= 4'd1;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd1;
        #(0*1s);
        addr0 <= 4'd10;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd6;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd2;
        #(0*1s);
        addr0 <= 4'd7;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd4;
        #(0*1s);
        web0 <= 1'b0;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        din0 <= 2'd0;
        #(0*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        addr0 <= 4'd2;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd1)) begin
            $error("Failed on action=196 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd1, dout0);
        end
        addr0 <= 4'd13;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=206 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd1;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=216 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd10;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd1)) begin
            $error("Failed on action=226 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd1, dout0);
        end
        addr0 <= 4'd7;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=236 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd14;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=246 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd11;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=256 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd15;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=266 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd8;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=276 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd4;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd0)) begin
            $error("Failed on action=286 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd0, dout0);
        end
        addr0 <= 4'd5;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=296 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd3;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=306 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd1)) begin
            $error("Failed on action=316 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd1, dout0);
        end
        addr0 <= 4'd9;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd3)) begin
            $error("Failed on action=326 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd3, dout0);
        end
        addr0 <= 4'd6;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd2)) begin
            $error("Failed on action=336 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd2, dout0);
        end
        addr0 <= 4'd12;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        #(1e-09*1s);
        clk0 <= 1'b1;
        #(0*1s);
        #(5e-09*1s);
        addr0 <= 4'd0;
        #(0*1s);
        web0 <= 1'b1;
        #(0*1s);
        clk0 <= 1'b0;
        #(0*1s);
        #(4e-09*1s);
        if (!(dout0 === 2'd1)) begin
            $error("Failed on action=346 checking port dout0 with traceback sram.py:116.  Expected %x, got %x.", 2'd1, dout0);
        end
        #20 $finish;
    end

endmodule

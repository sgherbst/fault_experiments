* Automatically generated file.
.include /home/sherbst/Code/OpenRAM/technology/scn4m_subm/models/nom/nmos.sp
.include /home/sherbst/Code/OpenRAM/technology/scn4m_subm/models/nom/pmos.sp
.include /home/sherbst/Code/fault_experiments/sram/build/temp/sram_2_16_scn4m_subm.sp
X0 din0[0] din0[1] addr0[0] addr0[1] addr0[2] addr0[3] csb0 web0 clk0 dout0[0] dout0[1] vdd gnd sram_2_16_scn4m_subm
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    Gs sw_p sw_n cur='V(sw_p, sw_n)*(0.999999999*V(ctl_p, ctl_n)+1e-09)'
.ends
X1 __din0[0]_v din0[0] __din0[0]_s 0 inout_sw_mod
V2 __din0[0]_v 0 DC 0 PWL(0 0 1e-07 0 1.002e-07 0 1.06e-07 0 1.062e-07 0 1.0999999999999999e-07 0 1.102e-07 3.3 1.1599999999999999e-07 3.3 1.162e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 0 1.46e-07 0 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 4.2000000000000027e-07 0)
V3 __din0[0]_s 0 DC 1 PWL(0 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 4.2000000000000027e-07 1)
X4 __din0[1]_v din0[1] __din0[1]_s 0 inout_sw_mod
V5 __din0[1]_v 0 DC 0 PWL(0 0 1e-07 0 1.002e-07 0 1.06e-07 0 1.062e-07 0 1.0999999999999999e-07 0 1.102e-07 3.3 1.1599999999999999e-07 3.3 1.162e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 0 1.46e-07 0 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 4.2000000000000027e-07 0)
V6 __din0[1]_s 0 DC 1 PWL(0 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 4.2000000000000027e-07 1)
X7 __addr0[0]_v addr0[0] __addr0[0]_s 0 inout_sw_mod
V8 __addr0[0]_v 0 DC 0 PWL(0 0 1e-07 0 1.002e-07 0 1.06e-07 0 1.062e-07 0 1.0999999999999999e-07 0 1.102e-07 0 1.1599999999999999e-07 0 1.162e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 0 2.7600000000000014e-07 0 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 0 2.9600000000000016e-07 0 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 0 3.160000000000002e-07 0 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 0 3.560000000000002e-07 0 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 0 3.6600000000000023e-07 0 3.6620000000000025e-07 0 3.700000000000002e-07 0 3.7020000000000023e-07 3.3 3.7600000000000024e-07 3.3 3.7620000000000026e-07 0 3.800000000000002e-07 0 3.8020000000000024e-07 0 3.8600000000000025e-07 0 3.8620000000000027e-07 0 3.9000000000000024e-07 0 3.9020000000000025e-07 0 3.9600000000000026e-07 0 3.962000000000003e-07 0 4.0000000000000025e-07 0 4.0020000000000026e-07 0 4.060000000000003e-07 0 4.062000000000003e-07 0 4.1000000000000026e-07 0 4.1020000000000027e-07 3.3 4.160000000000003e-07 3.3 4.162000000000003e-07 0 4.2000000000000027e-07 0)
V9 __addr0[0]_s 0 DC 1 PWL(0 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1 3.7020000000000023e-07 1 3.7600000000000024e-07 1 3.7620000000000026e-07 1 3.800000000000002e-07 1 3.8020000000000024e-07 1 3.8600000000000025e-07 1 3.8620000000000027e-07 1 3.9000000000000024e-07 1 3.9020000000000025e-07 1 3.9600000000000026e-07 1 3.962000000000003e-07 1 4.0000000000000025e-07 1 4.0020000000000026e-07 1 4.060000000000003e-07 1 4.062000000000003e-07 1 4.1000000000000026e-07 1 4.1020000000000027e-07 1 4.160000000000003e-07 1 4.162000000000003e-07 1 4.2000000000000027e-07 1)
X10 __addr0[1]_v addr0[1] __addr0[1]_s 0 inout_sw_mod
V11 __addr0[1]_v 0 DC 0 PWL(0 0 1e-07 0 1.002e-07 0 1.06e-07 0 1.062e-07 0 1.0999999999999999e-07 0 1.102e-07 0 1.1599999999999999e-07 0 1.162e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 0 1.46e-07 0 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 3.3 2.260000000000001e-07 3.3 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 0 3.360000000000002e-07 0 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 0 3.460000000000002e-07 0 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 0 3.560000000000002e-07 0 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 0 3.6600000000000023e-07 0 3.6620000000000025e-07 0 3.700000000000002e-07 0 3.7020000000000023e-07 0 3.7600000000000024e-07 0 3.7620000000000026e-07 0 3.800000000000002e-07 0 3.8020000000000024e-07 3.3 3.8600000000000025e-07 3.3 3.8620000000000027e-07 0 3.9000000000000024e-07 0 3.9020000000000025e-07 0 3.9600000000000026e-07 0 3.962000000000003e-07 0 4.0000000000000025e-07 0 4.0020000000000026e-07 0 4.060000000000003e-07 0 4.062000000000003e-07 0 4.1000000000000026e-07 0 4.1020000000000027e-07 0 4.160000000000003e-07 0 4.162000000000003e-07 0 4.2000000000000027e-07 0)
V12 __addr0[1]_s 0 DC 1 PWL(0 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1 3.7020000000000023e-07 1 3.7600000000000024e-07 1 3.7620000000000026e-07 1 3.800000000000002e-07 1 3.8020000000000024e-07 1 3.8600000000000025e-07 1 3.8620000000000027e-07 1 3.9000000000000024e-07 1 3.9020000000000025e-07 1 3.9600000000000026e-07 1 3.962000000000003e-07 1 4.0000000000000025e-07 1 4.0020000000000026e-07 1 4.060000000000003e-07 1 4.062000000000003e-07 1 4.1000000000000026e-07 1 4.1020000000000027e-07 1 4.160000000000003e-07 1 4.162000000000003e-07 1 4.2000000000000027e-07 1)
X13 __addr0[2]_v addr0[2] __addr0[2]_s 0 inout_sw_mod
V14 __addr0[2]_v 0 DC 0 PWL(0 0 1e-07 0 1.002e-07 3.3 1.06e-07 3.3 1.062e-07 0 1.0999999999999999e-07 0 1.102e-07 0 1.1599999999999999e-07 0 1.162e-07 0 1.2e-07 0 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 3.3 2.260000000000001e-07 3.3 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 0 2.6600000000000013e-07 0 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 0 2.7600000000000014e-07 0 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 0 3.160000000000002e-07 0 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 0 3.260000000000002e-07 0 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 0 3.460000000000002e-07 0 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 0 3.560000000000002e-07 0 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.700000000000002e-07 0 3.7020000000000023e-07 0 3.7600000000000024e-07 0 3.7620000000000026e-07 0 3.800000000000002e-07 0 3.8020000000000024e-07 3.3 3.8600000000000025e-07 3.3 3.8620000000000027e-07 0 3.9000000000000024e-07 0 3.9020000000000025e-07 0 3.9600000000000026e-07 0 3.962000000000003e-07 0 4.0000000000000025e-07 0 4.0020000000000026e-07 3.3 4.060000000000003e-07 3.3 4.062000000000003e-07 0 4.1000000000000026e-07 0 4.1020000000000027e-07 3.3 4.160000000000003e-07 3.3 4.162000000000003e-07 0 4.2000000000000027e-07 0)
V15 __addr0[2]_s 0 DC 1 PWL(0 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1 3.7020000000000023e-07 1 3.7600000000000024e-07 1 3.7620000000000026e-07 1 3.800000000000002e-07 1 3.8020000000000024e-07 1 3.8600000000000025e-07 1 3.8620000000000027e-07 1 3.9000000000000024e-07 1 3.9020000000000025e-07 1 3.9600000000000026e-07 1 3.962000000000003e-07 1 4.0000000000000025e-07 1 4.0020000000000026e-07 1 4.060000000000003e-07 1 4.062000000000003e-07 1 4.1000000000000026e-07 1 4.1020000000000027e-07 1 4.160000000000003e-07 1 4.162000000000003e-07 1 4.2000000000000027e-07 1)
X16 __addr0[3]_v addr0[3] __addr0[3]_s 0 inout_sw_mod
V17 __addr0[3]_v 0 DC 0 PWL(0 0 1e-07 0 1.002e-07 0 1.06e-07 0 1.062e-07 0 1.0999999999999999e-07 0 1.102e-07 0 1.1599999999999999e-07 0 1.162e-07 0 1.2e-07 0 1.2019999999999998e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.3e-07 0 1.302e-07 0 1.36e-07 0 1.362e-07 0 1.4e-07 0 1.402e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5000000000000002e-07 0 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 0 1.6000000000000003e-07 0 1.6020000000000002e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7000000000000004e-07 0 1.7020000000000003e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8000000000000005e-07 0 1.8020000000000004e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9000000000000006e-07 0 1.9020000000000005e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0000000000000007e-07 0 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 0 2.1000000000000008e-07 0 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 0 2.200000000000001e-07 0 2.2020000000000008e-07 3.3 2.260000000000001e-07 3.3 2.2620000000000008e-07 0 2.300000000000001e-07 0 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 0 2.400000000000001e-07 0 2.402000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 0 2.500000000000001e-07 0 2.502000000000001e-07 0 2.560000000000001e-07 0 2.5620000000000014e-07 0 2.600000000000001e-07 0 2.602000000000001e-07 0 2.6600000000000013e-07 0 2.6620000000000015e-07 0 2.700000000000001e-07 0 2.7020000000000013e-07 0 2.7600000000000014e-07 0 2.7620000000000016e-07 0 2.800000000000001e-07 0 2.8020000000000014e-07 0 2.8600000000000015e-07 0 2.8620000000000017e-07 0 2.9000000000000014e-07 0 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0000000000000015e-07 0 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.1000000000000016e-07 0 3.1020000000000017e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 0 3.2000000000000017e-07 0 3.202000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 0 3.300000000000002e-07 0 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.400000000000002e-07 0 3.402000000000002e-07 0 3.460000000000002e-07 0 3.4620000000000023e-07 0 3.500000000000002e-07 0 3.502000000000002e-07 0 3.560000000000002e-07 0 3.5620000000000024e-07 0 3.600000000000002e-07 0 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.700000000000002e-07 0 3.7020000000000023e-07 3.3 3.7600000000000024e-07 3.3 3.7620000000000026e-07 0 3.800000000000002e-07 0 3.8020000000000024e-07 0 3.8600000000000025e-07 0 3.8620000000000027e-07 0 3.9000000000000024e-07 0 3.9020000000000025e-07 3.3 3.9600000000000026e-07 3.3 3.962000000000003e-07 0 4.0000000000000025e-07 0 4.0020000000000026e-07 0 4.060000000000003e-07 0 4.062000000000003e-07 0 4.1000000000000026e-07 0 4.1020000000000027e-07 0 4.160000000000003e-07 0 4.162000000000003e-07 0 4.2000000000000027e-07 0)
V18 __addr0[3]_s 0 DC 1 PWL(0 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1 3.7020000000000023e-07 1 3.7600000000000024e-07 1 3.7620000000000026e-07 1 3.800000000000002e-07 1 3.8020000000000024e-07 1 3.8600000000000025e-07 1 3.8620000000000027e-07 1 3.9000000000000024e-07 1 3.9020000000000025e-07 1 3.9600000000000026e-07 1 3.962000000000003e-07 1 4.0000000000000025e-07 1 4.0020000000000026e-07 1 4.060000000000003e-07 1 4.062000000000003e-07 1 4.1000000000000026e-07 1 4.1020000000000027e-07 1 4.160000000000003e-07 1 4.162000000000003e-07 1 4.2000000000000027e-07 1)
X19 __csb0_v csb0 __csb0_s 0 inout_sw_mod
V20 __csb0_v 0 DC 0 PWL(0 0 4.2000000000000027e-07 0)
V21 __csb0_s 0 DC 1 PWL(0 1 4.2000000000000027e-07 1)
X22 __web0_v web0 __web0_s 0 inout_sw_mod
V23 __web0_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 1e-07 3.3 1.002e-07 0 1.06e-07 0 1.062e-07 3.3 1.0999999999999999e-07 3.3 1.102e-07 0 1.1599999999999999e-07 0 1.162e-07 3.3 1.2e-07 3.3 1.2019999999999998e-07 0 1.26e-07 0 1.2619999999999998e-07 3.3 1.3e-07 3.3 1.302e-07 0 1.36e-07 0 1.362e-07 3.3 1.4e-07 3.3 1.402e-07 0 1.46e-07 0 1.462e-07 3.3 1.5000000000000002e-07 3.3 1.502e-07 0 1.5600000000000002e-07 0 1.562e-07 3.3 1.6000000000000003e-07 3.3 1.6020000000000002e-07 0 1.6600000000000003e-07 0 1.6620000000000002e-07 3.3 1.7000000000000004e-07 3.3 1.7020000000000003e-07 0 1.7600000000000004e-07 0 1.7620000000000003e-07 3.3 1.8000000000000005e-07 3.3 1.8020000000000004e-07 0 1.8600000000000005e-07 0 1.8620000000000004e-07 3.3 1.9000000000000006e-07 3.3 1.9020000000000005e-07 0 1.9600000000000006e-07 0 1.9620000000000005e-07 3.3 2.0000000000000007e-07 3.3 2.0020000000000006e-07 0 2.0600000000000007e-07 0 2.0620000000000006e-07 3.3 2.1000000000000008e-07 3.3 2.1020000000000007e-07 0 2.1600000000000008e-07 0 2.1620000000000007e-07 3.3 2.200000000000001e-07 3.3 2.2020000000000008e-07 0 2.260000000000001e-07 0 2.2620000000000008e-07 3.3 2.300000000000001e-07 3.3 2.302000000000001e-07 0 2.360000000000001e-07 0 2.362000000000001e-07 3.3 2.400000000000001e-07 3.3 2.402000000000001e-07 0 2.460000000000001e-07 0 2.4620000000000013e-07 3.3 2.500000000000001e-07 3.3 2.502000000000001e-07 0 2.560000000000001e-07 0 2.5620000000000014e-07 3.3 2.600000000000001e-07 3.3 2.602000000000001e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 3.3 2.700000000000001e-07 3.3 2.7020000000000013e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 3.3 2.800000000000001e-07 3.3 2.8020000000000014e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 3.3 2.9000000000000014e-07 3.3 2.9020000000000015e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 3.3 3.0000000000000015e-07 3.3 3.0020000000000016e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 3.3 3.1000000000000016e-07 3.3 3.1020000000000017e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 3.3 3.2000000000000017e-07 3.3 3.202000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 3.3 3.300000000000002e-07 3.3 3.302000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 3.3 3.400000000000002e-07 3.3 3.402000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 3.3 3.500000000000002e-07 3.3 3.502000000000002e-07 3.3 3.560000000000002e-07 3.3 3.5620000000000024e-07 3.3 3.600000000000002e-07 3.3 3.602000000000002e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 3.3 3.700000000000002e-07 3.3 3.7020000000000023e-07 3.3 3.7600000000000024e-07 3.3 3.7620000000000026e-07 3.3 3.800000000000002e-07 3.3 3.8020000000000024e-07 3.3 3.8600000000000025e-07 3.3 3.8620000000000027e-07 3.3 3.9000000000000024e-07 3.3 3.9020000000000025e-07 3.3 3.9600000000000026e-07 3.3 3.962000000000003e-07 3.3 4.0000000000000025e-07 3.3 4.0020000000000026e-07 3.3 4.060000000000003e-07 3.3 4.062000000000003e-07 3.3 4.1000000000000026e-07 3.3 4.1020000000000027e-07 3.3 4.160000000000003e-07 3.3 4.162000000000003e-07 3.3 4.2000000000000027e-07 3.3)
V24 __web0_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 1e-07 1 1.002e-07 1 1.06e-07 1 1.062e-07 1 1.0999999999999999e-07 1 1.102e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2e-07 1 1.2019999999999998e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.3e-07 1 1.302e-07 1 1.36e-07 1 1.362e-07 1 1.4e-07 1 1.402e-07 1 1.46e-07 1 1.462e-07 1 1.5000000000000002e-07 1 1.502e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6000000000000003e-07 1 1.6020000000000002e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7000000000000004e-07 1 1.7020000000000003e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8000000000000005e-07 1 1.8020000000000004e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9000000000000006e-07 1 1.9020000000000005e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0000000000000007e-07 1 2.0020000000000006e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1000000000000008e-07 1 2.1020000000000007e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.200000000000001e-07 1 2.2020000000000008e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.300000000000001e-07 1 2.302000000000001e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.400000000000001e-07 1 2.402000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.500000000000001e-07 1 2.502000000000001e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.600000000000001e-07 1 2.602000000000001e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.700000000000001e-07 1 2.7020000000000013e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.800000000000001e-07 1 2.8020000000000014e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9000000000000014e-07 1 2.9020000000000015e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0000000000000015e-07 1 3.0020000000000016e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.1000000000000016e-07 1 3.1020000000000017e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.2000000000000017e-07 1 3.202000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.300000000000002e-07 1 3.302000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.400000000000002e-07 1 3.402000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.500000000000002e-07 1 3.502000000000002e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.600000000000002e-07 1 3.602000000000002e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.700000000000002e-07 1 3.7020000000000023e-07 1 3.7600000000000024e-07 1 3.7620000000000026e-07 1 3.800000000000002e-07 1 3.8020000000000024e-07 1 3.8600000000000025e-07 1 3.8620000000000027e-07 1 3.9000000000000024e-07 1 3.9020000000000025e-07 1 3.9600000000000026e-07 1 3.962000000000003e-07 1 4.0000000000000025e-07 1 4.0020000000000026e-07 1 4.060000000000003e-07 1 4.062000000000003e-07 1 4.1000000000000026e-07 1 4.1020000000000027e-07 1 4.160000000000003e-07 1 4.162000000000003e-07 1 4.2000000000000027e-07 1)
X25 __clk0_v clk0 __clk0_s 0 inout_sw_mod
V26 __clk0_v 0 DC 0 PWL(0 0 1.0099999999999999e-07 0 1.0119999999999999e-07 3.3 1.06e-07 3.3 1.062e-07 0 1.1099999999999999e-07 0 1.1119999999999999e-07 3.3 1.1599999999999999e-07 3.3 1.162e-07 0 1.2099999999999998e-07 0 1.2119999999999997e-07 3.3 1.26e-07 3.3 1.2619999999999998e-07 0 1.31e-07 0 1.3119999999999998e-07 3.3 1.36e-07 3.3 1.362e-07 0 1.41e-07 0 1.412e-07 3.3 1.46e-07 3.3 1.462e-07 0 1.5100000000000002e-07 0 1.512e-07 3.3 1.5600000000000002e-07 3.3 1.562e-07 0 1.6100000000000003e-07 0 1.6120000000000001e-07 3.3 1.6600000000000003e-07 3.3 1.6620000000000002e-07 0 1.7100000000000004e-07 0 1.7120000000000002e-07 3.3 1.7600000000000004e-07 3.3 1.7620000000000003e-07 0 1.8100000000000005e-07 0 1.8120000000000003e-07 3.3 1.8600000000000005e-07 3.3 1.8620000000000004e-07 0 1.9100000000000006e-07 0 1.9120000000000004e-07 3.3 1.9600000000000006e-07 3.3 1.9620000000000005e-07 0 2.0100000000000007e-07 0 2.0120000000000005e-07 3.3 2.0600000000000007e-07 3.3 2.0620000000000006e-07 0 2.1100000000000008e-07 0 2.1120000000000006e-07 3.3 2.1600000000000008e-07 3.3 2.1620000000000007e-07 0 2.2100000000000009e-07 0 2.2120000000000007e-07 3.3 2.260000000000001e-07 3.3 2.2620000000000008e-07 0 2.310000000000001e-07 0 2.3120000000000009e-07 3.3 2.360000000000001e-07 3.3 2.362000000000001e-07 0 2.410000000000001e-07 0 2.412000000000001e-07 3.3 2.460000000000001e-07 3.3 2.4620000000000013e-07 0 2.510000000000001e-07 0 2.5120000000000013e-07 3.3 2.560000000000001e-07 3.3 2.5620000000000014e-07 0 2.6100000000000013e-07 0 2.6120000000000014e-07 3.3 2.6600000000000013e-07 3.3 2.6620000000000015e-07 0 2.7100000000000014e-07 0 2.7120000000000015e-07 3.3 2.7600000000000014e-07 3.3 2.7620000000000016e-07 0 2.8100000000000015e-07 0 2.8120000000000016e-07 3.3 2.8600000000000015e-07 3.3 2.8620000000000017e-07 0 2.9100000000000016e-07 0 2.9120000000000017e-07 3.3 2.9600000000000016e-07 3.3 2.962000000000002e-07 0 3.0100000000000017e-07 0 3.012000000000002e-07 3.3 3.0600000000000017e-07 3.3 3.062000000000002e-07 0 3.110000000000002e-07 0 3.112000000000002e-07 3.3 3.160000000000002e-07 3.3 3.162000000000002e-07 0 3.210000000000002e-07 0 3.212000000000002e-07 3.3 3.260000000000002e-07 3.3 3.262000000000002e-07 0 3.310000000000002e-07 0 3.312000000000002e-07 3.3 3.360000000000002e-07 3.3 3.362000000000002e-07 0 3.410000000000002e-07 0 3.412000000000002e-07 3.3 3.460000000000002e-07 3.3 3.4620000000000023e-07 0 3.510000000000002e-07 0 3.5120000000000023e-07 3.3 3.560000000000002e-07 3.3 3.5620000000000024e-07 0 3.6100000000000023e-07 0 3.6120000000000024e-07 3.3 3.6600000000000023e-07 3.3 3.6620000000000025e-07 0 3.7100000000000024e-07 0 3.7120000000000025e-07 3.3 3.7600000000000024e-07 3.3 3.7620000000000026e-07 0 3.8100000000000025e-07 0 3.8120000000000026e-07 3.3 3.8600000000000025e-07 3.3 3.8620000000000027e-07 0 3.9100000000000026e-07 0 3.912000000000003e-07 3.3 3.9600000000000026e-07 3.3 3.962000000000003e-07 0 4.0100000000000027e-07 0 4.012000000000003e-07 3.3 4.060000000000003e-07 3.3 4.062000000000003e-07 0 4.110000000000003e-07 0 4.112000000000003e-07 3.3 4.160000000000003e-07 3.3 4.162000000000003e-07 0 4.2000000000000027e-07 0)
V27 __clk0_s 0 DC 1 PWL(0 1 1.0099999999999999e-07 1 1.0119999999999999e-07 1 1.06e-07 1 1.062e-07 1 1.1099999999999999e-07 1 1.1119999999999999e-07 1 1.1599999999999999e-07 1 1.162e-07 1 1.2099999999999998e-07 1 1.2119999999999997e-07 1 1.26e-07 1 1.2619999999999998e-07 1 1.31e-07 1 1.3119999999999998e-07 1 1.36e-07 1 1.362e-07 1 1.41e-07 1 1.412e-07 1 1.46e-07 1 1.462e-07 1 1.5100000000000002e-07 1 1.512e-07 1 1.5600000000000002e-07 1 1.562e-07 1 1.6100000000000003e-07 1 1.6120000000000001e-07 1 1.6600000000000003e-07 1 1.6620000000000002e-07 1 1.7100000000000004e-07 1 1.7120000000000002e-07 1 1.7600000000000004e-07 1 1.7620000000000003e-07 1 1.8100000000000005e-07 1 1.8120000000000003e-07 1 1.8600000000000005e-07 1 1.8620000000000004e-07 1 1.9100000000000006e-07 1 1.9120000000000004e-07 1 1.9600000000000006e-07 1 1.9620000000000005e-07 1 2.0100000000000007e-07 1 2.0120000000000005e-07 1 2.0600000000000007e-07 1 2.0620000000000006e-07 1 2.1100000000000008e-07 1 2.1120000000000006e-07 1 2.1600000000000008e-07 1 2.1620000000000007e-07 1 2.2100000000000009e-07 1 2.2120000000000007e-07 1 2.260000000000001e-07 1 2.2620000000000008e-07 1 2.310000000000001e-07 1 2.3120000000000009e-07 1 2.360000000000001e-07 1 2.362000000000001e-07 1 2.410000000000001e-07 1 2.412000000000001e-07 1 2.460000000000001e-07 1 2.4620000000000013e-07 1 2.510000000000001e-07 1 2.5120000000000013e-07 1 2.560000000000001e-07 1 2.5620000000000014e-07 1 2.6100000000000013e-07 1 2.6120000000000014e-07 1 2.6600000000000013e-07 1 2.6620000000000015e-07 1 2.7100000000000014e-07 1 2.7120000000000015e-07 1 2.7600000000000014e-07 1 2.7620000000000016e-07 1 2.8100000000000015e-07 1 2.8120000000000016e-07 1 2.8600000000000015e-07 1 2.8620000000000017e-07 1 2.9100000000000016e-07 1 2.9120000000000017e-07 1 2.9600000000000016e-07 1 2.962000000000002e-07 1 3.0100000000000017e-07 1 3.012000000000002e-07 1 3.0600000000000017e-07 1 3.062000000000002e-07 1 3.110000000000002e-07 1 3.112000000000002e-07 1 3.160000000000002e-07 1 3.162000000000002e-07 1 3.210000000000002e-07 1 3.212000000000002e-07 1 3.260000000000002e-07 1 3.262000000000002e-07 1 3.310000000000002e-07 1 3.312000000000002e-07 1 3.360000000000002e-07 1 3.362000000000002e-07 1 3.410000000000002e-07 1 3.412000000000002e-07 1 3.460000000000002e-07 1 3.4620000000000023e-07 1 3.510000000000002e-07 1 3.5120000000000023e-07 1 3.560000000000002e-07 1 3.5620000000000024e-07 1 3.6100000000000023e-07 1 3.6120000000000024e-07 1 3.6600000000000023e-07 1 3.6620000000000025e-07 1 3.7100000000000024e-07 1 3.7120000000000025e-07 1 3.7600000000000024e-07 1 3.7620000000000026e-07 1 3.8100000000000025e-07 1 3.8120000000000026e-07 1 3.8600000000000025e-07 1 3.8620000000000027e-07 1 3.9100000000000026e-07 1 3.912000000000003e-07 1 3.9600000000000026e-07 1 3.962000000000003e-07 1 4.0100000000000027e-07 1 4.012000000000003e-07 1 4.060000000000003e-07 1 4.062000000000003e-07 1 4.110000000000003e-07 1 4.112000000000003e-07 1 4.160000000000003e-07 1 4.162000000000003e-07 1 4.2000000000000027e-07 1)
X28 __vdd_v vdd __vdd_s 0 inout_sw_mod
V29 __vdd_v 0 DC 0 PWL(0 0 5e-08 0 5.02e-08 3.3 4.2000000000000027e-07 3.3)
V30 __vdd_s 0 DC 1 PWL(0 1 5e-08 1 5.02e-08 1 4.2000000000000027e-07 1)
X31 __gnd_v gnd __gnd_s 0 inout_sw_mod
V32 __gnd_v 0 DC 0 PWL(0 0 4.2000000000000027e-07 0)
V33 __gnd_s 0 DC 1 PWL(0 1 4.2000000000000027e-07 1)
.tran 4.2000000000000026e-10 4.2000000000000027e-07 uic
.control
run
set filetype=binary
write
exit
.endc
.probe V(dout0[1]) V(csb0) V(gnd) V(dout0[0]) V(addr0[0]) V(din0[0]) V(clk0) V(din0[1]) V(vdd) V(addr0[1]) V(web0) V(addr0[3]) V(addr0[2])
.end
